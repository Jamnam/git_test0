module a(
	input a,b;
	output c);
wire d;
wire e;

endmodule
